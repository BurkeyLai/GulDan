`timescale 1ns/10ps
`define CYCLE 10
/*
`include "DRAM.v"
*/

module top(
	/*
	your signal
	*/
);

/*
	DRAM DRAM_1 (
        .CK(clk),  
        .Q(Q),
        .RST(rst),
        .CSn(CSn),
        .WEn(WEn),
        .RASn(RASn),
        .CASn(CASn),
        .A(A),
        .D(D)
    );
*/

/*
	your code
*/


endmodule